library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- no entity
  -- no generics
  -- no ports


-- no architecture

  -- no signals

  -- no process
