library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity dummy is
  -- no generics
  -- no ports
end dummy;

-- no architecture

  -- no signals

  -- no process


