library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity dummy is
-- no generics
-- no ports
end dummy;

architecture behavioral of dummy is

-- no signals

begin

-- no process

end behavioral;